** sch_path: /foss/designs/DLL/2026/Cells/DLINE.sch
.subckt DLINE VSS VDD VIN VOUT
*.PININFO VOUT:O VIN:I VDD:B VSS:B
x7 net3 VIN VDD VSS sg13g2_dlygate4sd1_1
x7 net3 VIN VDD VSS sg13g2_dlygate4sd1_1
x9 net1 net VDD VSS sg13g2_inv_2
x9 net1 net VDD VSS sg13g2_inv_2
x9 net1 net VDD VSS sg13g2_inv_2
x9 net1 net VDD VSS sg13g2_inv_2
x1 net2 net VDD VSS sg13g2_inv_2
x1 net2 net VDD VSS sg13g2_inv_2
x1 net2 net VDD VSS sg13g2_inv_2
x1 net2 net VDD VSS sg13g2_inv_2
x1 net2 net VDD VSS sg13g2_inv_2
x1 net2 net VDD VSS sg13g2_inv_2
x1 net2 net VDD VSS sg13g2_inv_2
x1 net2 net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2
x2 VOUT net VDD VSS sg13g2_inv_2

* Library name: sg13g2_stdcell
* Cell name: sg13g2_dlygate4sd1_1
* View name: schematic
.subckt sg13g2_dlygate4sd1_1 X A VDD VSS
XP3 X net3 VDD VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=3.808e-13 as=3.808e-13 pd=2.92e-06 ps=2.92e-06 m=1
XP2 net3 net2 VDD VDD sg13_lv_pmos w=1.000u l=130.00n ng=1 ad=3.4e-13 as=3.4e-13 pd=2.68e-06 ps=2.68e-06 m=1
XP1 net2 net1 VDD VDD sg13_lv_pmos w=1.000u l=130.00n ng=1 ad=3.4e-13 as=3.4e-13 pd=2.68e-06 ps=2.68e-06 m=1
XP0 net1 A VDD VDD sg13_lv_pmos w=420.00n l=130.00n ng=1 ad=1.428e-13 as=1.428e-13 pd=1.52e-06 ps=1.52e-06 m=1
XN3 X net3 VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=2.516e-13 as=2.516e-13 pd=2.16e-06 ps=2.16e-06 m=1
XN2 net3 net2 VSS VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=1.428e-13 as=1.428e-13 pd=1.52e-06 ps=1.52e-06 m=1
XN1 net2 net1 VSS VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=1.428e-13 as=1.428e-13 pd=1.52e-06 ps=1.52e-06 m=1
XN0 net1 A VSS VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=1.428e-13 as=1.428e-13 pd=1.52e-06 ps=1.52e-06 m=1
.ends
* End of subcircuit definition.


* Library name: sg13g2_stdcell
* Cell name: sg13g2_inv_2
* View name: schematic
.subckt sg13g2_inv_2 Y A VDD VSS
MN1 Y A VSS VSS sg13_lv_nmos w=1.48u l=130.00n ng=2 ad=2.812e-13 as=5.032e-13 pd=2.24e-06 ps=4.32e-06 m=1
MP0 Y A VDD VDD sg13_lv_pmos w=2.24u l=130.00n ng=2 ad=4.256e-13 as=7.616e-13 pd=3e-06 ps=5.84e-06 m=1
.ends
* End of subcircuit definition.



.ends
