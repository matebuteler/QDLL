** sch_path: /foss/designs/DelayLine/xschem/QDLL.sch
.subckt QDLL VDD VSS IN1 OUT1 OUT2 IN2 CP
*.PININFO VDD:B VSS:B IN1:I IN2:I OUT1:O OUT2:O CP:B
x1 VDD OUT1 IN1 VSS CP TOP
x2 VDD OUT2 IN2 VSS CP TOP
x3 VSS OUT1 VDD OUT2 LATCH
.ends

* expanding   symbol:  Cells/TOP.sym # of pins=5
** sym_path: /foss/designs/DelayLine/xschem/Cells/TOP.sym
** sch_path: /foss/designs/DelayLine/xschem/Cells/TOP.sch
.subckt TOP VDD VOUT VIN VSS CP
*.PININFO VDD:B VOUT:O VIN:I VSS:B CP:B
x1 VSS VDD net1 VOUT DLine
x2 VDD VIN net1 CP VSS VCDL
x3 VDD VSS VIN net2 VOUT PD
x4 net2 CP VSS CP
.ends


* expanding   symbol:  Cells/LATCH.sym # of pins=4
** sym_path: /foss/designs/DelayLine/xschem/Cells/LATCH.sym
** sch_path: /foss/designs/DelayLine/xschem/Cells/LATCH.sch
.subckt LATCH VSS V1 VDD V2
*.PININFO VDD:B VSS:B V1:B V2:B
x1 V2 V1 VDD VSS sg13g2_inv_1
x2 V1 V2 VDD VSS sg13g2_inv_1
.ends


* expanding   symbol:  Cells/DLine.sym # of pins=4
** sym_path: /foss/designs/DelayLine/xschem/Cells/DLine.sym
** sch_path: /foss/designs/DelayLine/xschem/Cells/DLine.sch
.subckt DLine VSS VDD VIN VOUT
*.PININFO VOUT:O VIN:I VDD:B VSS:B
x7 net2 net1 VDD VSS sg13g2_dlygate4sd1_1
x1 net2 net1 VDD VSS sg13g2_dlygate4sd1_1
x2 net3 net2 VDD VSS sg13g2_inv_4
x3 net4 net3 VDD VSS sg13g2_inv_8
x4 VOUT net4 VDD VSS sg13g2_inv_16
x5 net1 net7 VDD VSS sg13g2_dlygate4sd1_1
x6 net7 net6 VDD VSS sg13g2_dlygate4sd1_1
x8 net6 net5 VDD VSS sg13g2_dlygate4sd1_1
x9 net5 VIN VDD VSS sg13g2_dlygate4sd1_1
.ends


* expanding   symbol:  Cells/VCDL.sym # of pins=5
** sym_path: /foss/designs/DelayLine/xschem/Cells/VCDL.sym
** sch_path: /foss/designs/DelayLine/xschem/Cells/VCDL.sch
.subckt VCDL VDD VIN VOUT VCONT VSS
*.PININFO VDD:B VSS:B VIN:I VCONT:I VOUT:O
XM1 VOUT VIN net3 VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM2 net3 VCONT VSS VSS sg13_lv_nmos w=3.5u l=0.18u ng=1 m=1
XM3 net1 VCONT VSS VSS sg13_lv_nmos w=2u l=0.25u ng=1 m=1
XM4 VOUT VIN net2 VDD sg13_lv_pmos w=4.46u l=0.13u ng=1 m=1
Xq net2 net1 VDD VDD sg13_lv_pmos w=2.24u l=0.13u ng=1 m=1
XM6 net1 net1 VDD VDD sg13_lv_pmos w=2.24u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  Cells/PD.sym # of pins=5
** sym_path: /foss/designs/DelayLine/xschem/Cells/PD.sym
** sch_path: /foss/designs/DelayLine/xschem/Cells/PD.sch
.subckt PD VDD VSS PDIN1 PDOUT PDIN2
*.PININFO VDD:B VSS:B PDOUT:O PDIN1:I PDIN2:I
x1 PDOUT PDIN1 PDIN2 VDD VSS sg13g2_xor2_1
.ends


* expanding   symbol:  Cells/CP.sym # of pins=3
** sym_path: /foss/designs/DelayLine/xschem/Cells/CP.sym
** sch_path: /foss/designs/DelayLine/xschem/Cells/CP.sch
.subckt CP CPIN CPOUT VSS
*.PININFO VSS:B CPIN:I CPOUT:O
XC1 CPOUT VSS cap_cmim w=20e-6 l=20e-6 m=1
x1 net1 CPIN RES
x2 CPOUT net1 RES
XC2 CPOUT VSS cap_cmim w=20e-6 l=20e-6 m=1
XC3 CPOUT VSS cap_cmim w=20e-6 l=20e-6 m=1
.ends


* expanding   symbol:  Cells/RES.sym # of pins=2
** sym_path: /foss/designs/DelayLine/xschem/Cells/RES.sym
** sch_path: /foss/designs/DelayLine/xschem/Cells/RES.sch
.subckt RES ROUT RIN
*.PININFO RIN:I ROUT:O
XR1 net1 RIN sub! rppd w=1e-6 l=10e-6 m=1 b=0
XR3 net2 net1 sub! rppd w=1e-6 l=10e-6 m=1 b=0
XR4 net3 net2 sub! rppd w=1e-6 l=10e-6 m=1 b=0
XR5 ROUT net3 sub! rppd w=1e-6 l=10e-6 m=1 b=0
.ends

