** CACE Template: Phase Detector Characterization
** sch_path: tb_pd.sch

.param vdd_val = CACE{vdd}
.param temp_val = CACE{temperature}

** Include PDK models
.lib CACE{PDK_ROOT}/CACE{PDK}/libs.tech/ngspice/models/cornerMOSlv.lib mos_CACE{corner}
.lib CACE{PDK_ROOT}/CACE{PDK}/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib CACE{PDK_ROOT}/CACE{PDK}/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.include CACE{PDK_ROOT}/CACE{PDK}/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

** Include DUT (Phase Detector subcircuit)
.include "CACE{DUT_path}"

** Temperature
.temp CACE{temperature}

** Power supplies
Vdd VDD GND CACE{vdd}
Vss VSS GND 0

** Reference clock (fixed)
Vref CK_REF GND PULSE(0 CACE{vdd} 0 10p 10p 1n 2n)

** Input clock with variable phase (sweep phase)
Vin CK_IN GND PULSE(0 CACE{vdd} 0.5n 10p 10p 1n 2n)

** DUT instance - Phase Detector
XPD CK_IN UP CK_REF DN CACE{DUT_name}

** Charge pump load
Ccp VC GND 1p

** Analysis
.tran 1p 20n

** Measure average voltages to calculate gain
.meas tran vup_avg AVG v(UP) FROM=10n TO=20n
.meas tran vdn_avg AVG v(DN) FROM=10n TO=20n
.meas tran pd_gain PARAM='(vup_avg-vdn_avg)/0.785'

** Output results
.control
run
set filetype=ascii
echo $&pd_gain > CACE{simpath}/CACE{filename}_CACE{N}.data
.endc

.end