** CACE Template: Power Consumption Measurement
** sch_path: tb_power.sch

.param vdd_val = CACE{vdd}
.param temp_val = CACE{temperature}
.param fin_val = CACE{fin}

** Include PDK models
.lib CACE{PDK_ROOT}/CACE{PDK}/libs.tech/ngspice/models/cornerMOSlv.lib mos_CACE{corner}
.lib CACE{PDK_ROOT}/CACE{PDK}/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib CACE{PDK_ROOT}/CACE{PDK}/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.include CACE{PDK_ROOT}/CACE{PDK}/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

** Include DUT
.include "CACE{DUT_path}"

** Temperature
.temp CACE{temperature}

** Power supplies with current measurement
Vdd VDD GND CACE{vdd}
Vss VSS GND 0

** Clock inputs at specified frequency
.param period_ns = '1000/CACE{fin}'
Vin1 IN1 GND PULSE(0 CACE{vdd} 0 10p 10p 'period_ns/2*1n' 'period_ns*1n')
Vin2 IN2 GND PULSE(0 CACE{vdd} 'period_ns/4*1n' 10p 10p 'period_ns/2*1n' 'period_ns*1n')

** Control voltage set to 0.6 V as a mid-range "typical" operating point for the DLL
** This value was chosen based on nominal PVT characterization; sweep externally if needed
Vcont CP GND 0.6

** DUT instance - using QDLL
XDUT VDD VSS IN1 IN2 OUT1 OUT2 CP QDLL

** Load capacitors
Cload1 OUT1 GND 100f
Cload2 OUT2 GND 100f

** Analysis - static then dynamic
.tran 10p 200n

** Measurements
.meas tran idd_static AVG i(Vdd) FROM=0n TO=10n
.meas tran idd_dynamic AVG i(Vdd) FROM=100n TO=200n

** Output results (convert to uA and mA)
.control
run
let idd_static_ua = abs(idd_static) * 1e6
let idd_dynamic_ma = abs(idd_dynamic) * 1e3
set filetype=ascii
echo $&idd_static_ua $&idd_dynamic_ma > CACE{simpath}/CACE{filename}_CACE{N}.data
.endc

.end