-- sch_path: /foss/designs/DLL/2026/Cells/RES.sch
entity RES is
port(
  ROUT : out std_logic ;
  RIN :  in std_logic
);
end RES ;

architecture arch_RES of RES is


signal sub! : std_logic ;
signal VSS : std_logic ;
signal net1 : std_logic ;
signal net2 : std_logic ;
signal net3 : std_logic ;
begin
end arch_RES ;

