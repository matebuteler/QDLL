** sch_path: /foss/designs/UNIC-CASS-Aug25/sch/delay_variable_line/variable_delay_line.sch
**.subckt variable_delay_line VDD VSS VCONT VOUT VIN
*.iopin VSS
*.iopin VDD
*.ipin VIN
*.opin VOUT
*.ipin VCONT
x1 VDD VIN va VCONT VSS delay_variable
x2 VDD VSS va VOUT large_delay_vto1p1
**.ends

* expanding   symbol:  /foss/designs/UNIC-CASS-Aug25/sch/delay_variable/delay_variable.sym # of pins=5
** sym_path: /foss/designs/UNIC-CASS-Aug25/sch/delay_variable/delay_variable.sym
** sch_path: /foss/designs/UNIC-CASS-Aug25/sch/delay_variable/delay_variable.sch
.subckt delay_variable VDD_D VIN_D VOUT_D VCONT_D VSS_D
*.iopin VDD_D
*.opin VOUT_D
*.ipin VCONT_D
*.ipin VIN_D
*.iopin VSS_D
XM3 net3 VCONT_D VSS_D VSS_D sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM5 net2 VCONT_D VSS_D VSS_D sg13_lv_nmos w=2u l=2u ng=1 m=1
XM4 net3 net3 VDD_D VDD_D sg13_lv_pmos w=2.24u l=0.13u ng=1 m=1
XM6 net1 net3 VDD_D VDD_D sg13_lv_pmos w=4u l=2u ng=1 m=1
XM7 VOUT_D VIN_D net1 VDD_D sg13_lv_pmos w=4u l=2u ng=4 m=1
XM8 VOUT_D VIN_D net2 VSS_D sg13_lv_nmos w=5u l=3u ng=1 m=1
.ends


* expanding   symbol:  /foss/designs/UNIC-CASS-Aug25/sch/large_delay_vto1p1/large_delay_vto1p1.sym # of pins=4
** sym_path: /foss/designs/UNIC-CASS-Aug25/sch/large_delay_vto1p1/large_delay_vto1p1.sym
** sch_path: /foss/designs/UNIC-CASS-Aug25/sch/large_delay_vto1p1/large_delay_vto1p1.sch
.subckt large_delay_vto1p1 VCC VSS VIN VOUT
*.iopin VIN
*.iopin VOUT
*.iopin VCC
*.iopin VSS
x1 VIN VCC VSS net1 sg13g2_dlygate4sd1_1
x2 VIN VCC VSS net1 sg13g2_dlygate4sd1_1
x3 VIN VCC VSS net1 sg13g2_dlygate4sd1_1
x4 VIN VCC VSS net1 sg13g2_dlygate4sd1_1
x5 net1 VCC VSS VOUT sg13g2_dlygate4sd3_1
.ends

.end
