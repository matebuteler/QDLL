* Extracted by KLayout with SG13G2 LVS runset on : 24/01/2026 08:59

.SUBCKT DLYGATES2 VSS A|VIN VOUT|X VDD
M$1 \$3 A|VIN VSS VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.1428p
+ PS=1.52u PD=1.1u
M$2 VSS \$3 \$4 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.1428p PS=1.1u
+ PD=1.52u
M$3 VSS \$4 \$5 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1405p AD=0.2373p PS=1.15u
+ PD=1.97u
M$4 VSS \$5 VOUT|X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1405p AD=0.2516p
+ PS=1.15u PD=2.16u
M$5 \$10 \$9 VSS VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1405p
+ PS=1.97u PD=1.15u
M$6 VSS \$10 VOUT|X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1405p AD=0.2516p
+ PS=1.15u PD=2.16u
M$7 \$8 A|VIN VSS VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.1428p
+ PS=1.52u PD=1.1u
M$8 VSS \$8 \$9 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.1428p PS=1.1u
+ PD=1.52u
M$9 VDD A|VIN \$3 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.2931p AD=0.1428p
+ PS=1.65u PD=1.52u
M$10 VDD \$3 \$4 VDD sg13_lv_pmos L=0.13u W=1u AS=0.2931p AD=0.37p PS=1.65u
+ PD=2.74u
M$11 \$5 \$4 VDD VDD sg13_lv_pmos L=0.13u W=1u AS=0.565p AD=0.2245p PS=3.13u
+ PD=1.53u
M$12 VDD \$5 VOUT|X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2245p AD=0.3808p
+ PS=1.53u PD=2.92u
M$13 VDD A|VIN \$8 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.2931p AD=0.1428p
+ PS=1.65u PD=1.52u
M$14 VDD \$8 \$9 VDD sg13_lv_pmos L=0.13u W=1u AS=0.2931p AD=0.37p PS=1.65u
+ PD=2.74u
M$15 VDD \$9 \$10 VDD sg13_lv_pmos L=0.13u W=1u AS=0.2245p AD=0.565p PS=1.53u
+ PD=3.13u
M$16 VDD \$10 VOUT|X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2245p AD=0.3808p
+ PS=1.53u PD=2.92u
.ENDS DLYGATES2
