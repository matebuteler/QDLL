** sch_path: /foss/designs/DLL/2026/Cells/TOP.sch
**.subckt TOP VDD VOUT VIN VCONT VSS CPOUT PD2
*.iopin VDD
*.opin VOUT
*.ipin VCONT
*.ipin VIN
*.iopin VSS
*.ipin PD2
*.opin CPOUT
x1 VSS VDD net1 VOUT DLine
x2 VDD VIN net1 VCONT VSS VCDL
x3 VDD VSS VIN net2 PD2 PD
x4 net2 CPOUT VSS CP
**.ends

* expanding   symbol:  /foss/designs/DLL/2026/Cells/DLine.sym # of pins=4
** sym_path: /foss/designs/DLL/2026/Cells/DLine.sym
** sch_path: /foss/designs/DLL/2026/Cells/DLine.sch
.subckt DLine VSS VDD VIN VOUT
*.opin VOUT
*.ipin VIN
*.iopin VDD
*.iopin VSS
x7[1] net3_1 VIN VDD VSS sg13g2_dlygate4sd1_1
x7[0] net3_0 VIN VDD VSS sg13g2_dlygate4sd1_1
x9[3] net1_3 net3_1 VDD VSS sg13g2_inv_2
x9[2] net1_2 net3_0 VDD VSS sg13g2_inv_2
x9[1] net1_1 net3_1 VDD VSS sg13g2_inv_2
x9[0] net1_0 net3_0 VDD VSS sg13g2_inv_2
x1[7] net2_7 net1_3 VDD VSS sg13g2_inv_2
x1[6] net2_6 net1_2 VDD VSS sg13g2_inv_2
x1[5] net2_5 net1_1 VDD VSS sg13g2_inv_2
x1[4] net2_4 net1_0 VDD VSS sg13g2_inv_2
x1[3] net2_3 net1_3 VDD VSS sg13g2_inv_2
x1[2] net2_2 net1_2 VDD VSS sg13g2_inv_2
x1[1] net2_1 net1_1 VDD VSS sg13g2_inv_2
x1[0] net2_0 net1_0 VDD VSS sg13g2_inv_2
x2[15] VOUT net2_7 VDD VSS sg13g2_inv_2
x2[14] VOUT net2_6 VDD VSS sg13g2_inv_2
x2[13] VOUT net2_5 VDD VSS sg13g2_inv_2
x2[12] VOUT net2_4 VDD VSS sg13g2_inv_2
x2[11] VOUT net2_3 VDD VSS sg13g2_inv_2
x2[10] VOUT net2_2 VDD VSS sg13g2_inv_2
x2[9] VOUT net2_1 VDD VSS sg13g2_inv_2
x2[8] VOUT net2_0 VDD VSS sg13g2_inv_2
x2[7] VOUT net2_7 VDD VSS sg13g2_inv_2
x2[6] VOUT net2_6 VDD VSS sg13g2_inv_2
x2[5] VOUT net2_5 VDD VSS sg13g2_inv_2
x2[4] VOUT net2_4 VDD VSS sg13g2_inv_2
x2[3] VOUT net2_3 VDD VSS sg13g2_inv_2
x2[2] VOUT net2_2 VDD VSS sg13g2_inv_2
x2[1] VOUT net2_1 VDD VSS sg13g2_inv_2
x2[0] VOUT net2_0 VDD VSS sg13g2_inv_2
.ends


* expanding   symbol:  /foss/designs/DLL/2026/Cells/VCDL.sym # of pins=5
** sym_path: /foss/designs/DLL/2026/Cells/VCDL.sym
** sch_path: /foss/designs/DLL/2026/Cells/VCDL.sch
.subckt VCDL VDD VIN VOUT VCONT VSS
*.iopin VDD
*.iopin VSS
*.ipin VIN
*.ipin VCONT
*.opin VOUT
XM1 VOUT VIN net3 VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM2 net3 VCONT VSS VSS sg13_lv_nmos w=2u l=0.16u ng=1 m=1
XM3 net1 VCONT VSS VSS sg13_lv_nmos w=2u l=0.25u ng=1 m=1
XM4 VOUT VIN net2 VDD sg13_lv_pmos w=4.46u l=0.13u ng=1 m=1
XM5 net2 net1 VDD VDD sg13_lv_pmos w=1.5u l=0.16u ng=1 m=1
XM6 net1 net1 VDD VDD sg13_lv_pmos w=2.24u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /foss/designs/DLL/2026/Cells/PD.sym # of pins=5
** sym_path: /foss/designs/DLL/2026/Cells/PD.sym
** sch_path: /foss/designs/DLL/2026/Cells/PD.sch
.subckt PD VDD VSS PDIN1 PDOUT PDIN2
*.iopin VDD
*.iopin VSS
*.opin PDOUT
*.ipin PDIN1
*.ipin PDIN2
x1 PDOUT PDIN1 PDIN2 VDD VSS sg13g2_xor2_1
.ends


* expanding   symbol:  /foss/designs/DLL/2026/Cells/CP.sym # of pins=3
** sym_path: /foss/designs/DLL/2026/Cells/CP.sym
** sch_path: /foss/designs/DLL/2026/Cells/CP.sch
.subckt CP CPIN CPOUT VSS
*.iopin VSS
*.ipin CPIN
*.opin CPOUT
XC1 CPOUT VSS cap_cmim w=20e-6 l=20e-6 m=1
x1 net1 CPIN RES
x2 CPOUT net1 RES
.ends


* expanding   symbol:  /foss/designs/DLL/2026/Cells/RES.sym # of pins=2
** sym_path: /foss/designs/DLL/2026/Cells/RES.sym
** sch_path: /foss/designs/DLL/2026/Cells/RES.sch
.subckt RES ROUT RIN
*.ipin RIN
*.opin ROUT
XR1 net1 RIN sub! rppd w=1e-6 l=10e-6 m=1 b=0
XR3 net2 net1 sub! rppd w=1e-6 l=10e-6 m=1 b=0
XR4 net3 net2 sub! rppd w=1e-6 l=10e-6 m=1 b=0
XR5 ROUT net3 sub! rppd w=1e-6 l=10e-6 m=1 b=0
.ends




* Library name: sg13g2_stdcell
* Cell name: sg13g2_xor2_1
* View name: schematic
.subckt sg13g2_xor2_1 X A B VDD VSS
MN0 net1 A VSS VSS sg13_lv_nmos w=550.00n l=130.00n ng=1 ad=1.87e-13 as=1.87e-13 pd=1.78e-06 ps=1.78e-06 m=1
MN4 X B net3 VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=2.516e-13 as=2.516e-13 pd=2.16e-06 ps=2.16e-06 m=1
MN6 X net1 VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=2.516e-13 as=2.516e-13 pd=2.16e-06 ps=2.16e-06 m=1
MN8 net3 A VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=2.516e-13 as=2.516e-13 pd=2.16e-06 ps=2.16e-06 m=1
MN9 net1 B VSS VSS sg13_lv_nmos w=550.00n l=130.00n ng=1 ad=1.87e-13 as=1.87e-13 pd=1.78e-06 ps=1.78e-06 m=1
MP1 net6 A VDD VDD sg13_lv_pmos w=1.000u l=130.00n ng=1 ad=3.4e-13 as=3.4e-13 pd=2.68e-06 ps=2.68e-06 m=1
MP2 net1 B net6 VDD sg13_lv_pmos w=1.000u l=130.00n ng=1 ad=3.4e-13 as=3.4e-13 pd=2.68e-06 ps=2.68e-06 m=1
MP3 net5 A VDD VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=3.808e-13 as=3.808e-13 pd=2.92e-06 ps=2.92e-06 m=1
MP5 net5 B VDD VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=3.808e-13 as=3.808e-13 pd=2.92e-06 ps=2.92e-06 m=1
MP7 X net1 net5 VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=3.808e-13 as=3.808e-13 pd=2.92e-06 ps=2.92e-06 m=1
.ends
* End of subcircuit definition.

* Library name: sg13g2_stdcell
* Cell name: sg13g2_dlygate4sd1_1
* View name: schematic
.subckt sg13g2_dlygate4sd1_1 X A VDD VSS
MP3 X net3 VDD VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=3.808e-13 as=3.808e-13 pd=2.92e-06 ps=2.92e-06 m=1
MP2 net3 net2 VDD VDD sg13_lv_pmos w=1.000u l=130.00n ng=1 ad=3.4e-13 as=3.4e-13 pd=2.68e-06 ps=2.68e-06 m=1
MP1 net2 net1 VDD VDD sg13_lv_pmos w=1.000u l=130.00n ng=1 ad=3.4e-13 as=3.4e-13 pd=2.68e-06 ps=2.68e-06 m=1
MP0 net1 A VDD VDD sg13_lv_pmos w=420.00n l=130.00n ng=1 ad=1.428e-13 as=1.428e-13 pd=1.52e-06 ps=1.52e-06 m=1
MN3 X net3 VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=2.516e-13 as=2.516e-13 pd=2.16e-06 ps=2.16e-06 m=1
MN2 net3 net2 VSS VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=1.428e-13 as=1.428e-13 pd=1.52e-06 ps=1.52e-06 m=1
MN1 net2 net1 VSS VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=1.428e-13 as=1.428e-13 pd=1.52e-06 ps=1.52e-06 m=1
MN0 net1 A VSS VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=1.428e-13 as=1.428e-13 pd=1.52e-06 ps=1.52e-06 m=1
.ends
* End of subcircuit definition.


* Library name: sg13g2_stdcell
* Cell name: sg13g2_inv_2
* View name: schematic
.subckt sg13g2_inv_2 Y A VDD VSS
MN1 Y A VSS VSS sg13_lv_nmos w=1.48u l=130.00n ng=2 ad=2.812e-13 as=5.032e-13 pd=2.24e-06 ps=4.32e-06 m=1
MP0 Y A VDD VDD sg13_lv_pmos w=2.24u l=130.00n ng=2 ad=4.256e-13 as=7.616e-13 pd=3e-06 ps=5.84e-06 m=1
.ends
* End of subcircuit definition.



.end
