** sch_path: /foss/designs/DLL/2026/example/nor3_res.sch
**.subckt nor3_res VOUT VA VB VC
*.iopin VOUT
*.iopin VA
*.iopin VB
*.iopin VC
x1 net1 VA VB VC VDD VSS sg13g2_nor3_1
XR1 net1 VOUT sub! rppd w=0.5e-6 l=0.5e-6 m=1 b=0
**.ends

* Library name: sg13g2_stdcell
* Cell name: sg13g2_nor3_1
* View name: schematic
.subckt sg13g2_nor3_1 Y A B C VDD VSS
MP3 Y C net2 VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=3.808e-13 as=3.808e-13 pd=2.92e-06 ps=2.92e-06 m=1
MP0 net2 B net3 VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=3.808e-13 as=3.808e-13 pd=2.92e-06 ps=2.92e-06 m=1
MP2 net3 A VDD VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=3.808e-13 as=3.808e-13 pd=2.92e-06 ps=2.92e-06 m=1
MN4 Y A VSS VSS sg13_lv_nmos w=770.00n l=130.00n ng=1 ad=2.618e-13 as=2.618e-13 pd=2.22e-06 ps=2.22e-06 m=1
MN1 Y B VSS VSS sg13_lv_nmos w=770.00n l=130.00n ng=1 ad=2.618e-13 as=2.618e-13 pd=2.22e-06 ps=2.22e-06 m=1
MN5 Y C VSS VSS sg13_lv_nmos w=770.00n l=130.00n ng=1 ad=2.618e-13 as=2.618e-13 pd=2.22e-06 ps=2.22e-06 m=1
.ends
* End of subcircuit definition.



.end
