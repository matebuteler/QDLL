** sch_path: /foss/designs/DelayLine/cace/templates/tb_pd.sch
**.subckt tb_pd
Vdd VDD GND CACE{vdd}
Vref CK_REF GND PULSE(0 CACE{vdd} 0 10p 10p 1n 2n)
Vin CK_IN GND PULSE(0 CACE{vdd} 0.5n 10p 10p 1n 2n)
x1 VDD GND CK_IN net1 CK_REF PD
**** begin user architecture code

.param vdd_val=1.2

.param vdd_val = CACE{vdd}
.param temp_val = CACE{temperature}

** Include PDK models
.lib CACE{PDK_ROOT}/CACE{PDK}/libs.tech/ngspice/models/cornerMOSlv.lib mos_CACE{corner}
.lib CACE{PDK_ROOT}/CACE{PDK}/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib CACE{PDK_ROOT}/CACE{PDK}/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.include CACE{PDK_ROOT}/CACE{PDK}/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

** Include DUT (Phase Detector subcircuit)
.include CACE{DUT_path}

** Temperature
.temp CACE{temperature}

** Analysis
.tran 1p 20n

** Measure average voltages to calculate gain
.meas tran vup_avg AVG v(UP) FROM=10n TO=20n
.meas tran vdn_avg AVG v(DN) FROM=10n TO=20n
.meas tran pd_gain PARAM='(vup_avg-vdn_avg)/0.785'

** Output results
.control
run
set filetype=ascii
echo $&pd_gain > CACE{simpath}/CACE{filename}_CACE{N}.data
.endc

.end

**** end user architecture code
**.ends

* expanding   symbol:  Cells/PD.sym # of pins=5
** sym_path: /foss/designs/DelayLine/xschem/Cells/PD.sym
** sch_path: /foss/designs/DelayLine/xschem/Cells/PD.sch
.subckt PD VDD VSS PDIN1 PDOUT PDIN2
*.iopin VDD
*.iopin VSS
*.opin PDOUT
*.ipin PDIN1
*.ipin PDIN2
x1 PDOUT PDIN1 PDIN2 VDD VSS sg13g2_xor2_1
.ends

.GLOBAL GND
.end
