** sch_path: /foss/designs/DLL/2026/Cells/VCDL.sch
.subckt VCDL VDD VIN VOUT VCONT VSS
*.PININFO VDD:B VSS:B VIN:I VCONT:I VOUT:O
M1 VOUT VIN net3 VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
M2 net3 VCONT VSS VSS sg13_lv_nmos w=3.5u l=0.16u ng=1 m=1
M3 net1 VCONT VSS VSS sg13_lv_nmos w=2u l=0.25u ng=1 m=1
M4 VOUT VIN net2 VDD sg13_lv_pmos w=4.46u l=0.13u ng=1 m=1
M5 net2 net1 VDD VDD sg13_lv_pmos w=2.8u l=0.16u ng=1 m=1
M6 net1 net1 VDD VDD sg13_lv_pmos w=2.24u l=0.13u ng=1 m=1
.ends
