** sch_path: /foss/designs/DLL/2026/Cells/INV4.sch
**.subckt INV4 VSS VDD VOUT VIN
*.ipin VIN
*.iopin VDD
*.iopin VSS
*.opin VOUT
x9 VOUT VIN VDD VSS sg13g2_inv_2
x2 VOUT VIN VDD VSS sg13g2_inv_2
x3 VOUT VIN VDD VSS sg13g2_inv_2
x4 VOUT VIN VDD VSS sg13g2_inv_2
**.ends


* Library name: sg13g2_stdcell
* Cell name: sg13g2_inv_2
* View name: schematic
.subckt sg13g2_inv_2 Y A VDD VSS
MN1 Y A VSS VSS sg13_lv_nmos w=1.48u l=130.00n ng=2 ad=2.812e-13 as=5.032e-13 pd=2.24e-06 ps=4.32e-06 m=1
MP0 Y A VDD VDD sg13_lv_pmos w=2.24u l=130.00n ng=2 ad=4.256e-13 as=7.616e-13 pd=3e-06 ps=5.84e-06 m=1
.ends
* End of subcircuit definition.



.end
