* Extracted by KLayout with SG13G2 LVS runset on : 24/01/2026 10:06

.SUBCKT INV16 VSS A|VOUT VIN|Y VDD
M$1 VSS A|VOUT VIN|Y VSS sg13_lv_nmos L=0.13u W=11.84u AS=2.3606p AD=2.3606p
+ PS=18.96u PD=18.96u
M$17 VDD A|VOUT VIN|Y VDD sg13_lv_pmos L=0.13u W=17.92u AS=3.5728p AD=3.6288p
+ PS=25.42u PD=25.52u
.ENDS INV16
